library verilog;
use verilog.vl_types.all;
entity testTcircuit is
end testTcircuit;
